// Dump of memory (4 banks in parallel)
localparam [DQ_BITS : 0] in_mem [ 0 : 8191][0 : 3]  = '{
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hffff, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hffff, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hffff, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hffff } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'hf800, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'h07e0, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hf800, 16'h001f, 16'h001f, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'hffff, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hffff, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hffff, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h07e0, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h001f, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hf800, 16'hf800, 16'h001f, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'hf800, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'h07e0, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hf800 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'h07e0 } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hffff } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'h001f } ,
  '{16'h001f, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hf800, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'h07e0, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hffff, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'h001f, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'h07e0, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'h001f, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'h001f, 16'hf800, 16'hxxxx, 16'hxxxx } ,
  '{16'hffff, 16'hffff, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hf800, 16'h07e0, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } ,
  '{16'hxxxx, 16'hxxxx, 16'hxxxx, 16'hxxxx } };
